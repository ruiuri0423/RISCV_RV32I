module LSU #(

)(

);

endmodule